// This is just a stub to satisfy the IP flow 
module pxi_ii_wizard_v1_0_1_top(
	output wiz
); 

endmodule


